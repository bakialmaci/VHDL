--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:49:09 12/01/2018
-- Design Name:   
-- Module Name:   D:/Xilinx/three_eight_decoder/ted_tb.vhd
-- Project Name:  three_eight_decoder
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: three_eight_decoder
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY ted_tb IS
END ted_tb;
 
ARCHITECTURE behavior OF ted_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT three_eight_decoder
    PORT(
         x : IN  std_logic;
         y : IN  std_logic;
         z : IN  std_logic;
         d : OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal x : std_logic := '0';
   signal y : std_logic := '0';
   signal z : std_logic := '0';

 	--Outputs
   signal d : std_logic_vector(7 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
--   constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: three_eight_decoder PORT MAP (
          x => x,
          y => y,
          z => z,
          d => d
        );

   -- Clock process definitions
--   <clock>_process :process
--   begin
--		<clock> <= '0';
--		wait for <clock>_period/2;
--		<clock> <= '1';
--		wait for <clock>_period/2;
--   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      x <= '0';
		y <= '0';
		z <= '0';
      wait for 100 ns;	
      x <= '0';
		y <= '0';
		z <= '1';
      wait for 100 ns;
      x <= '0';
		y <= '1';
		z <= '0';
      wait for 100 ns;
      x <= '0';
		y <= '1';
		z <= '1';
      wait for 100 ns;
      x <= '1';
		y <= '0';
		z <= '0';
      wait for 100 ns;
      x <= '1';
		y <= '0';
		z <= '1';
      wait for 100 ns;
      x <= '1';
		y <= '1';
		z <= '0';
      wait for 100 ns;
      x <= '1';
		y <= '1';
		z <= '1';
      wait;
   end process;

END;
